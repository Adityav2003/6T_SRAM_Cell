magic
tech sky130A
timestamp 1712003917
<< nwell >>
rect -35 200 70 310
rect 325 200 430 310
rect -35 100 130 200
rect 265 100 430 200
<< nmos >>
rect 40 -110 55 -10
rect 340 -110 355 -10
rect 80 -165 160 -150
rect 235 -165 315 -150
<< pmos >>
rect 40 120 55 180
rect 340 120 355 180
<< ndiff >>
rect -35 -35 40 -10
rect -35 -90 -20 -35
rect 20 -90 40 -35
rect -35 -110 40 -90
rect 55 -20 130 -10
rect 55 -65 75 -20
rect 100 -65 130 -20
rect 55 -110 130 -65
rect 265 -20 340 -10
rect 265 -65 295 -20
rect 320 -65 340 -20
rect 265 -110 340 -65
rect 355 -35 430 -10
rect 355 -90 375 -35
rect 415 -90 430 -35
rect 355 -110 430 -90
rect 80 -150 160 -110
rect 235 -150 315 -110
rect 80 -185 160 -165
rect 80 -205 100 -185
rect 140 -205 160 -185
rect 80 -210 160 -205
rect 235 -185 315 -165
rect 235 -205 255 -185
rect 295 -205 315 -185
rect 235 -210 315 -205
<< pdiff >>
rect -15 165 40 180
rect -15 135 0 165
rect 20 135 40 165
rect -15 120 40 135
rect 55 170 110 180
rect 55 130 75 170
rect 100 130 110 170
rect 55 120 110 130
rect 285 170 340 180
rect 285 130 295 170
rect 320 130 340 170
rect 285 120 340 130
rect 355 165 410 180
rect 355 135 375 165
rect 395 135 410 165
rect 355 120 410 135
<< ndiffc >>
rect -20 -90 20 -35
rect 75 -65 100 -20
rect 295 -65 320 -20
rect 375 -90 415 -35
rect 100 -205 140 -185
rect 255 -205 295 -185
<< pdiffc >>
rect 0 135 20 165
rect 75 130 100 170
rect 295 130 320 170
rect 375 135 395 165
<< psubdiff >>
rect -30 -155 30 -145
rect -30 -180 -15 -155
rect 15 -180 30 -155
rect 365 -155 425 -145
rect -30 -190 30 -180
rect 365 -180 380 -155
rect 410 -180 425 -155
rect 365 -190 425 -180
<< nsubdiff >>
rect -15 275 35 290
rect -15 225 -5 275
rect 25 225 35 275
rect -15 210 35 225
rect 360 275 410 290
rect 360 225 370 275
rect 400 225 410 275
rect 360 210 410 225
<< psubdiffcont >>
rect -15 -180 15 -155
rect 380 -180 410 -155
<< nsubdiffcont >>
rect -5 225 25 275
rect 370 225 400 275
<< poly >>
rect 40 180 55 195
rect 340 180 355 195
rect 40 35 55 120
rect 340 90 355 120
rect 80 85 355 90
rect 80 65 90 85
rect 110 65 355 85
rect 80 60 355 65
rect 40 30 315 35
rect 40 10 285 30
rect 305 10 315 30
rect 40 5 315 10
rect 40 -10 55 5
rect 340 -10 355 60
rect 40 -125 55 -110
rect 340 -125 355 -110
rect 65 -165 80 -150
rect 160 -165 235 -150
rect 315 -165 330 -150
rect 180 -185 215 -165
rect 180 -210 185 -185
rect 210 -210 215 -185
rect 180 -220 215 -210
<< polycont >>
rect 90 65 110 85
rect 285 10 305 30
rect 185 -210 210 -185
<< locali >>
rect -15 285 35 290
rect 360 285 410 290
rect -15 280 410 285
rect -15 275 180 280
rect -15 225 -5 275
rect 25 250 180 275
rect 215 275 410 280
rect 215 250 370 275
rect 25 245 370 250
rect 25 225 35 245
rect -15 210 35 225
rect 360 225 370 245
rect 400 225 410 275
rect 360 210 410 225
rect -10 165 30 210
rect -10 135 0 165
rect 20 135 30 165
rect -10 125 30 135
rect 65 170 110 180
rect 65 130 75 170
rect 100 130 110 170
rect 65 85 110 130
rect 65 65 90 85
rect 65 -20 110 65
rect -30 -35 30 -25
rect -30 -90 -20 -35
rect 20 -90 30 -35
rect 65 -65 75 -20
rect 100 -65 110 -20
rect 65 -75 110 -65
rect 285 170 330 180
rect 285 130 295 170
rect 320 130 330 170
rect 285 30 330 130
rect 365 165 405 210
rect 365 135 375 165
rect 395 135 405 165
rect 365 125 405 135
rect 305 10 330 30
rect 285 -20 330 10
rect 285 -65 295 -20
rect 320 -65 330 -20
rect 285 -75 330 -65
rect 365 -35 425 -25
rect -30 -155 30 -90
rect -30 -180 -15 -155
rect 15 -180 30 -155
rect 365 -90 375 -35
rect 415 -90 425 -35
rect 365 -155 425 -90
rect -30 -190 30 -180
rect 90 -185 150 -175
rect 245 -185 305 -175
rect 90 -205 100 -185
rect 140 -205 150 -185
rect 90 -235 150 -205
rect 90 -265 105 -235
rect 135 -265 150 -235
rect 175 -210 185 -185
rect 210 -210 220 -185
rect 175 -235 220 -210
rect 175 -260 185 -235
rect 210 -260 220 -235
rect 175 -265 220 -260
rect 245 -205 255 -185
rect 295 -205 305 -185
rect 365 -180 380 -155
rect 410 -180 425 -155
rect 365 -190 425 -180
rect 245 -235 305 -205
rect 245 -265 260 -235
rect 290 -265 305 -235
<< viali >>
rect 180 250 215 280
rect -10 -175 10 -155
rect 105 -265 135 -235
rect 185 -260 210 -235
rect 385 -175 405 -155
rect 260 -265 290 -235
<< metal1 >>
rect 145 280 250 360
rect 145 250 180 280
rect 215 250 250 280
rect 145 230 250 250
rect -35 -155 35 -145
rect -35 -175 -10 -155
rect 10 -175 35 -155
rect -35 -235 35 -175
rect 360 -155 430 -145
rect 360 -175 385 -155
rect 405 -175 430 -155
rect 85 -235 155 -230
rect 85 -265 105 -235
rect 135 -265 155 -235
rect 85 -305 155 -265
rect 175 -235 220 -230
rect 175 -260 185 -235
rect 210 -260 220 -235
rect 175 -335 220 -260
rect 240 -235 310 -230
rect 360 -235 430 -175
rect 240 -265 260 -235
rect 290 -265 310 -235
rect 240 -305 310 -265
<< labels >>
rlabel metal1 195 325 195 325 1 vdd
rlabel metal1 390 -215 390 -215 1 gnd
rlabel metal1 -15 -215 -15 -215 1 gnd
rlabel metal1 195 -315 195 -315 1 wl
rlabel metal1 115 -290 115 -290 1 bl
rlabel metal1 275 -290 275 -290 1 blb
<< end >>
